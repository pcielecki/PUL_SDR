--
--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 
--
--   To use any of the example code shown below, uncomment the lines and modify as necessary
--

library IEEE;
use IEEE.STD_LOGIC_1164.all;

package sin_lut_pkg is

type sin_lut_array is array (511 downto 0) of integer range 0 to (2**16-1);

constant lut_array : sin_lut_array := (32768,
33170,
33572,
33974,
34375,
34777,
35178,
35579,
35979,
36379,
36779,
37177,
37575,
37973,
38369,
38765,
39160,
39554,
39947,
40339,
40729,
41119,
41507,
41894,
42279,
42663,
43046,
43427,
43807,
44184,
44560,
44935,
45307,
45678,
46046,
46413,
46777,
47140,
47500,
47858,
48214,
48567,
48919,
49267,
49613,
49957,
50298,
50636,
50972,
51305,
51635,
51963,
52287,
52609,
52927,
53243,
53555,
53864,
54170,
54473,
54773,
55069,
55362,
55652,
55938,
56220,
56499,
56775,
57047,
57315,
57579,
57840,
58097,
58350,
58600,
58845,
59087,
59324,
59558,
59787,
60013,
60234,
60451,
60664,
60873,
61078,
61278,
61474,
61666,
61853,
62036,
62215,
62389,
62559,
62724,
62885,
63041,
63192,
63339,
63482,
63620,
63753,
63881,
64005,
64124,
64238,
64348,
64453,
64553,
64648,
64739,
64825,
64905,
64981,
65053,
65119,
65180,
65237,
65289,
65335,
65377,
65414,
65446,
65473,
65496,
65513,
65525,
65533,
65535,
65533,
65525,
65513,
65496,
65473,
65446,
65414,
65377,
65335,
65289,
65237,
65180,
65119,
65053,
64981,
64905,
64825,
64739,
64648,
64553,
64453,
64348,
64238,
64124,
64005,
63881,
63753,
63620,
63482,
63339,
63192,
63041,
62885,
62724,
62559,
62389,
62215,
62036,
61853,
61666,
61474,
61278,
61078,
60873,
60664,
60451,
60234,
60013,
59787,
59558,
59324,
59087,
58845,
58600,
58350,
58097,
57840,
57579,
57315,
57047,
56775,
56499,
56220,
55938,
55652,
55362,
55069,
54773,
54473,
54170,
53864,
53555,
53243,
52927,
52609,
52287,
51963,
51635,
51305,
50972,
50636,
50298,
49957,
49613,
49267,
48919,
48567,
48214,
47858,
47500,
47140,
46777,
46413,
46046,
45678,
45307,
44935,
44560,
44184,
43807,
43427,
43046,
42663,
42279,
41894,
41507,
41119,
40729,
40339,
39947,
39554,
39160,
38765,
38369,
37973,
37575,
37177,
36779,
36379,
35979,
35579,
35178,
34777,
34375,
33974,
33572,
33170,
32768,
32365,
31963,
31561,
31160,
30758,
30357,
29956,
29556,
29156,
28756,
28358,
27960,
27562,
27166,
26770,
26375,
25981,
25588,
25196,
24806,
24416,
24028,
23641,
23256,
22872,
22489,
22108,
21728,
21351,
20975,
20600,
20228,
19857,
19489,
19122,
18758,
18395,
18035,
17677,
17321,
16968,
16616,
16268,
15922,
15578,
15237,
14899,
14563,
14230,
13900,
13572,
13248,
12926,
12608,
12292,
11980,
11671,
11365,
11062,
10762,
10466,
10173,
9883,
9597,
9315,
9036,
8760,
8488,
8220,
7956,
7695,
7438,
7185,
6935,
6690,
6448,
6211,
5977,
5748,
5522,
5301,
5084,
4871,
4662,
4457,
4257,
4061,
3869,
3682,
3499,
3320,
3146,
2976,
2811,
2650,
2494,
2343,
2196,
2053,
1915,
1782,
1654,
1530,
1411,
1297,
1187,
1082,
982,
887,
796,
710,
630,
554,
482,
416,
355,
298,
246,
200,
158,
121,
89,
62,
39,
22,
10,
2,
0,
2,
10,
22,
39,
62,
89,
121,
158,
200,
246,
298,
355,
416,
482,
554,
630,
710,
796,
887,
982,
1082,
1187,
1297,
1411,
1530,
1654,
1782,
1915,
2053,
2196,
2343,
2494,
2650,
2811,
2976,
3146,
3320,
3499,
3682,
3869,
4061,
4257,
4457,
4662,
4871,
5084,
5301,
5522,
5748,
5977,
6211,
6448,
6690,
6935,
7185,
7438,
7695,
7956,
8220,
8488,
8760,
9036,
9315,
9597,
9883,
10173,
10466,
10762,
11062,
11365,
11671,
11980,
12292,
12608,
12926,
13248,
13572,
13900,
14230,
14563,
14899,
15237,
15578,
15922,
16268,
16616,
16968,
17321,
17677,
18035,
18395,
18758,
19122,
19489,
19857,
20228,
20600,
20975,
21351,
21728,
22108,
22489,
22872,
23256,
23641,
24028,
24416,
24806,
25196,
25588,
25981,
26375,
26770,
27166,
27562,
27960,
28358,
28756,
29156,
29556,
29956,
30357,
30758,
31160,
31561,
31963,
32365);

end sin_lut_pkg;

package body sin_lut_pkg is

---- Example 1
--  function <function_name>  (signal <signal_name> : in <type_declaration>  ) return <type_declaration> is
--    variable <variable_name>     : <type_declaration>;
--  begin
--    <variable_name> := <signal_name> xor <signal_name>;
--    return <variable_name>; 
--  end <function_name>;

---- Example 2
--  function <function_name>  (signal <signal_name> : in <type_declaration>;
--                         signal <signal_name>   : in <type_declaration>  ) return <type_declaration> is
--  begin
--    if (<signal_name> = '1') then
--      return <signal_name>;
--    else
--      return 'Z';
--    end if;
--  end <function_name>;

---- Procedure Example
--  procedure <procedure_name>  (<type_declaration> <constant_name>  : in <type_declaration>) is
--    
--  begin
--    
--  end <procedure_name>;
 
end sin_lut_pkg;

--
--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 
--
--   To use any of the example code shown below, uncomment the lines and modify as necessary
--

library IEEE;
use IEEE.STD_LOGIC_1164.all;

package sin_lut_pkg is

type sin_lut_array is array (0 to 1389) of integer range 0 to (2**16-1);

constant lut_array : sin_lut_array := (32768,
32916,
33064,
33212,
33360,
33508,
33656,
33804,
33952,
34100,
34248,
34396,
34544,
34692,
34840,
34988,
35135,
35283,
35431,
35578,
35726,
35873,
36021,
36168,
36315,
36463,
36610,
36757,
36904,
37051,
37197,
37344,
37491,
37637,
37784,
37930,
38076,
38222,
38368,
38514,
38660,
38806,
38951,
39097,
39242,
39387,
39532,
39677,
39822,
39966,
40111,
40255,
40399,
40543,
40687,
40830,
40974,
41117,
41260,
41403,
41546,
41689,
41831,
41973,
42115,
42257,
42399,
42540,
42682,
42823,
42964,
43104,
43245,
43385,
43525,
43665,
43804,
43944,
44083,
44222,
44360,
44499,
44637,
44775,
44913,
45050,
45187,
45324,
45461,
45597,
45733,
45869,
46005,
46140,
46275,
46410,
46545,
46679,
46813,
46947,
47080,
47213,
47346,
47478,
47611,
47743,
47874,
48005,
48136,
48267,
48397,
48527,
48657,
48786,
48916,
49044,
49173,
49301,
49428,
49556,
49683,
49809,
49936,
50062,
50187,
50313,
50438,
50562,
50686,
50810,
50934,
51057,
51179,
51302,
51424,
51545,
51667,
51787,
51908,
52028,
52147,
52267,
52385,
52504,
52622,
52740,
52857,
52974,
53090,
53206,
53322,
53437,
53551,
53666,
53780,
53893,
54006,
54119,
54231,
54342,
54454,
54565,
54675,
54785,
54894,
55003,
55112,
55220,
55328,
55435,
55542,
55648,
55754,
55859,
55964,
56068,
56172,
56275,
56378,
56481,
56583,
56684,
56785,
56886,
56986,
57085,
57184,
57283,
57381,
57479,
57576,
57672,
57768,
57864,
57959,
58053,
58147,
58240,
58333,
58426,
58518,
58609,
58700,
58790,
58880,
58969,
59058,
59146,
59233,
59320,
59407,
59493,
59578,
59663,
59748,
59831,
59915,
59997,
60079,
60161,
60242,
60322,
60402,
60482,
60560,
60638,
60716,
60793,
60870,
60945,
61021,
61095,
61170,
61243,
61316,
61389,
61460,
61532,
61602,
61672,
61742,
61811,
61879,
61947,
62014,
62080,
62146,
62212,
62276,
62340,
62404,
62467,
62529,
62591,
62652,
62712,
62772,
62831,
62890,
62948,
63005,
63062,
63118,
63174,
63228,
63283,
63336,
63389,
63442,
63494,
63545,
63595,
63645,
63694,
63743,
63791,
63838,
63885,
63931,
63977,
64022,
64066,
64109,
64152,
64194,
64236,
64277,
64317,
64357,
64396,
64434,
64472,
64509,
64546,
64581,
64617,
64651,
64685,
64718,
64751,
64783,
64814,
64844,
64874,
64904,
64932,
64960,
64987,
65014,
65040,
65065,
65090,
65114,
65137,
65160,
65182,
65203,
65224,
65244,
65263,
65282,
65300,
65318,
65334,
65350,
65366,
65380,
65394,
65408,
65420,
65433,
65444,
65455,
65465,
65474,
65483,
65491,
65498,
65505,
65511,
65516,
65521,
65525,
65528,
65531,
65533,
65534,
65535,
65535,
65534,
65533,
65531,
65528,
65525,
65521,
65516,
65511,
65505,
65498,
65491,
65483,
65474,
65465,
65455,
65444,
65433,
65420,
65408,
65394,
65380,
65366,
65350,
65334,
65318,
65300,
65282,
65263,
65244,
65224,
65203,
65182,
65160,
65137,
65114,
65090,
65065,
65040,
65014,
64987,
64960,
64932,
64904,
64874,
64844,
64814,
64783,
64751,
64718,
64685,
64651,
64617,
64581,
64546,
64509,
64472,
64434,
64396,
64357,
64317,
64277,
64236,
64194,
64152,
64109,
64066,
64022,
63977,
63931,
63885,
63838,
63791,
63743,
63694,
63645,
63595,
63545,
63494,
63442,
63389,
63336,
63283,
63228,
63174,
63118,
63062,
63005,
62948,
62890,
62831,
62772,
62712,
62652,
62591,
62529,
62467,
62404,
62340,
62276,
62212,
62146,
62080,
62014,
61947,
61879,
61811,
61742,
61672,
61602,
61532,
61460,
61389,
61316,
61243,
61170,
61095,
61021,
60945,
60870,
60793,
60716,
60638,
60560,
60482,
60402,
60322,
60242,
60161,
60079,
59997,
59915,
59831,
59748,
59663,
59578,
59493,
59407,
59320,
59233,
59146,
59058,
58969,
58880,
58790,
58700,
58609,
58518,
58426,
58333,
58240,
58147,
58053,
57959,
57864,
57768,
57672,
57576,
57479,
57381,
57283,
57184,
57085,
56986,
56886,
56785,
56684,
56583,
56481,
56378,
56275,
56172,
56068,
55964,
55859,
55754,
55648,
55542,
55435,
55328,
55220,
55112,
55003,
54894,
54785,
54675,
54565,
54454,
54342,
54231,
54119,
54006,
53893,
53780,
53666,
53551,
53437,
53322,
53206,
53090,
52974,
52857,
52740,
52622,
52504,
52385,
52267,
52147,
52028,
51908,
51787,
51667,
51545,
51424,
51302,
51179,
51057,
50934,
50810,
50686,
50562,
50438,
50313,
50187,
50062,
49936,
49809,
49683,
49556,
49428,
49301,
49173,
49044,
48916,
48786,
48657,
48527,
48397,
48267,
48136,
48005,
47874,
47743,
47611,
47478,
47346,
47213,
47080,
46947,
46813,
46679,
46545,
46410,
46275,
46140,
46005,
45869,
45733,
45597,
45461,
45324,
45187,
45050,
44913,
44775,
44637,
44499,
44360,
44222,
44083,
43944,
43804,
43665,
43525,
43385,
43245,
43104,
42964,
42823,
42682,
42540,
42399,
42257,
42115,
41973,
41831,
41689,
41546,
41403,
41260,
41117,
40974,
40830,
40687,
40543,
40399,
40255,
40111,
39966,
39822,
39677,
39532,
39387,
39242,
39097,
38951,
38806,
38660,
38514,
38368,
38222,
38076,
37930,
37784,
37637,
37491,
37344,
37197,
37051,
36904,
36757,
36610,
36463,
36315,
36168,
36021,
35873,
35726,
35578,
35431,
35283,
35135,
34988,
34840,
34692,
34544,
34396,
34248,
34100,
33952,
33804,
33656,
33508,
33360,
33212,
33064,
32916,
32768,
32619,
32471,
32323,
32175,
32027,
31879,
31731,
31583,
31435,
31287,
31139,
30991,
30843,
30695,
30547,
30400,
30252,
30104,
29957,
29809,
29662,
29514,
29367,
29220,
29072,
28925,
28778,
28631,
28484,
28338,
28191,
28044,
27898,
27751,
27605,
27459,
27313,
27167,
27021,
26875,
26729,
26584,
26438,
26293,
26148,
26003,
25858,
25713,
25569,
25424,
25280,
25136,
24992,
24848,
24705,
24561,
24418,
24275,
24132,
23989,
23846,
23704,
23562,
23420,
23278,
23136,
22995,
22853,
22712,
22571,
22431,
22290,
22150,
22010,
21870,
21731,
21591,
21452,
21313,
21175,
21036,
20898,
20760,
20622,
20485,
20348,
20211,
20074,
19938,
19802,
19666,
19530,
19395,
19260,
19125,
18990,
18856,
18722,
18588,
18455,
18322,
18189,
18057,
17924,
17792,
17661,
17530,
17399,
17268,
17138,
17008,
16878,
16749,
16619,
16491,
16362,
16234,
16107,
15979,
15852,
15726,
15599,
15473,
15348,
15222,
15097,
14973,
14849,
14725,
14601,
14478,
14356,
14233,
14111,
13990,
13868,
13748,
13627,
13507,
13388,
13268,
13150,
13031,
12913,
12795,
12678,
12561,
12445,
12329,
12213,
12098,
11984,
11869,
11755,
11642,
11529,
11416,
11304,
11193,
11081,
10970,
10860,
10750,
10641,
10532,
10423,
10315,
10207,
10100,
9993,
9887,
9781,
9676,
9571,
9467,
9363,
9260,
9157,
9054,
8952,
8851,
8750,
8649,
8549,
8450,
8351,
8252,
8154,
8056,
7959,
7863,
7767,
7671,
7576,
7482,
7388,
7295,
7202,
7109,
7017,
6926,
6835,
6745,
6655,
6566,
6477,
6389,
6302,
6215,
6128,
6042,
5957,
5872,
5787,
5704,
5620,
5538,
5456,
5374,
5293,
5213,
5133,
5053,
4975,
4897,
4819,
4742,
4665,
4590,
4514,
4440,
4365,
4292,
4219,
4146,
4075,
4003,
3933,
3863,
3793,
3724,
3656,
3588,
3521,
3455,
3389,
3323,
3259,
3195,
3131,
3068,
3006,
2944,
2883,
2823,
2763,
2704,
2645,
2587,
2530,
2473,
2417,
2361,
2307,
2252,
2199,
2146,
2093,
2041,
1990,
1940,
1890,
1841,
1792,
1744,
1697,
1650,
1604,
1558,
1513,
1469,
1426,
1383,
1341,
1299,
1258,
1218,
1178,
1139,
1101,
1063,
1026,
989,
954,
918,
884,
850,
817,
784,
752,
721,
691,
661,
631,
603,
575,
548,
521,
495,
470,
445,
421,
398,
375,
353,
332,
311,
291,
272,
253,
235,
217,
201,
185,
169,
155,
141,
127,
115,
102,
91,
80,
70,
61,
52,
44,
37,
30,
24,
19,
14,
10,
7,
4,
2,
1,
0,
0,
1,
2,
4,
7,
10,
14,
19,
24,
30,
37,
44,
52,
61,
70,
80,
91,
102,
115,
127,
141,
155,
169,
185,
201,
217,
235,
253,
272,
291,
311,
332,
353,
375,
398,
421,
445,
470,
495,
521,
548,
575,
603,
631,
661,
691,
721,
752,
784,
817,
850,
884,
918,
954,
989,
1026,
1063,
1101,
1139,
1178,
1218,
1258,
1299,
1341,
1383,
1426,
1469,
1513,
1558,
1604,
1650,
1697,
1744,
1792,
1841,
1890,
1940,
1990,
2041,
2093,
2146,
2199,
2252,
2307,
2361,
2417,
2473,
2530,
2587,
2645,
2704,
2763,
2823,
2883,
2944,
3006,
3068,
3131,
3195,
3259,
3323,
3389,
3455,
3521,
3588,
3656,
3724,
3793,
3863,
3933,
4003,
4075,
4146,
4219,
4292,
4365,
4440,
4514,
4590,
4665,
4742,
4819,
4897,
4975,
5053,
5133,
5213,
5293,
5374,
5456,
5538,
5620,
5704,
5787,
5872,
5957,
6042,
6128,
6215,
6302,
6389,
6477,
6566,
6655,
6745,
6835,
6926,
7017,
7109,
7202,
7295,
7388,
7482,
7576,
7671,
7767,
7863,
7959,
8056,
8154,
8252,
8351,
8450,
8549,
8649,
8750,
8851,
8952,
9054,
9157,
9260,
9363,
9467,
9571,
9676,
9781,
9887,
9993,
10100,
10207,
10315,
10423,
10532,
10641,
10750,
10860,
10970,
11081,
11193,
11304,
11416,
11529,
11642,
11755,
11869,
11984,
12098,
12213,
12329,
12445,
12561,
12678,
12795,
12913,
13031,
13150,
13268,
13388,
13507,
13627,
13748,
13868,
13990,
14111,
14233,
14356,
14478,
14601,
14725,
14849,
14973,
15097,
15222,
15348,
15473,
15599,
15726,
15852,
15979,
16107,
16234,
16362,
16491,
16619,
16749,
16878,
17008,
17138,
17268,
17399,
17530,
17661,
17792,
17924,
18057,
18189,
18322,
18455,
18588,
18722,
18856,
18990,
19125,
19260,
19395,
19530,
19666,
19802,
19938,
20074,
20211,
20348,
20485,
20622,
20760,
20898,
21036,
21175,
21313,
21452,
21591,
21731,
21870,
22010,
22150,
22290,
22431,
22571,
22712,
22853,
22995,
23136,
23278,
23420,
23562,
23704,
23846,
23989,
24132,
24275,
24418,
24561,
24705,
24848,
24992,
25136,
25280,
25424,
25569,
25713,
25858,
26003,
26148,
26293,
26438,
26584,
26729,
26875,
27021,
27167,
27313,
27459,
27605,
27751,
27898,
28044,
28191,
28338,
28484,
28631,
28778,
28925,
29072,
29220,
29367,
29514,
29662,
29809,
29957,
30104,
30252,
30400,
30547,
30695,
30843,
30991,
31139,
31287,
31435,
31583,
31731,
31879,
32027,
32175,
32323,
32471,
32619);

end sin_lut_pkg;

package body sin_lut_pkg is

---- Example 1
--  function <function_name>  (signal <signal_name> : in <type_declaration>  ) return <type_declaration> is
--    variable <variable_name>     : <type_declaration>;
--  begin
--    <variable_name> := <signal_name> xor <signal_name>;
--    return <variable_name>; 
--  end <function_name>;

---- Example 2
--  function <function_name>  (signal <signal_name> : in <type_declaration>;
--                         signal <signal_name>   : in <type_declaration>  ) return <type_declaration> is
--  begin
--    if (<signal_name> = '1') then
--      return <signal_name>;
--    else
--      return 'Z';
--    end if;
--  end <function_name>;

---- Procedure Example
--  procedure <procedure_name>  (<type_declaration> <constant_name>  : in <type_declaration>) is
--    
--  begin
--    
--  end <procedure_name>;
 
end sin_lut_pkg;

--
--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 
--
--   To use any of the example code shown below, uncomment the lines and modify as necessary
--

library IEEE;
use IEEE.STD_LOGIC_1164.all;

package sin_lut_pkg is

type sin_lut_array is array (0 to 1389) of integer range (- 2**15) to (2**15-1);

constant lut_array : sin_lut_array := (
0,
147,
295,
443,
591,
740,
888,
1036,
1184,
1332,
1480,
1628,
1776,
1923,
2071,
2219,
2367,
2515,
2662,
2810,
2957,
3105,
3252,
3400,
3547,
3694,
3841,
3988,
4135,
4282,
4429,
4576,
4722,
4869,
5015,
5162,
5308,
5454,
5600,
5746,
5892,
6037,
6183,
6328,
6473,
6619,
6764,
6908,
7053,
7198,
7342,
7486,
7631,
7775,
7918,
8062,
8205,
8349,
8492,
8635,
8778,
8920,
9063,
9205,
9347,
9489,
9631,
9772,
9913,
10054,
10195,
10336,
10476,
10617,
10757,
10896,
11036,
11175,
11315,
11453,
11592,
11730,
11869,
12007,
12144,
12282,
12419,
12556,
12693,
12829,
12965,
13101,
13237,
13372,
13507,
13642,
13776,
13911,
14045,
14178,
14312,
14445,
14578,
14710,
14842,
14974,
15106,
15237,
15368,
15499,
15629,
15759,
15889,
16018,
16147,
16276,
16404,
16532,
16660,
16788,
16915,
17041,
17168,
17294,
17419,
17544,
17669,
17794,
17918,
18042,
18165,
18289,
18411,
18534,
18656,
18777,
18898,
19019,
19140,
19260,
19379,
19498,
19617,
19736,
19854,
19971,
20089,
20205,
20322,
20438,
20553,
20668,
20783,
20898,
21011,
21125,
21238,
21350,
21463,
21574,
21686,
21796,
21907,
22017,
22126,
22235,
22344,
22452,
22559,
22667,
22773,
22880,
22985,
23091,
23196,
23300,
23404,
23507,
23610,
23713,
23815,
23916,
24017,
24118,
24218,
24317,
24416,
24515,
24613,
24710,
24807,
24904,
25000,
25095,
25190,
25285,
25379,
25472,
25565,
25658,
25749,
25841,
25932,
26022,
26112,
26201,
26290,
26378,
26465,
26552,
26639,
26725,
26810,
26895,
26979,
27063,
27146,
27229,
27311,
27393,
27474,
27554,
27634,
27713,
27792,
27870,
27948,
28025,
28101,
28177,
28253,
28327,
28402,
28475,
28548,
28621,
28692,
28764,
28834,
28904,
28974,
29043,
29111,
29179,
29246,
29312,
29378,
29443,
29508,
29572,
29636,
29699,
29761,
29823,
29884,
29944,
30004,
30063,
30122,
30180,
30237,
30294,
30350,
30406,
30460,
30515,
30568,
30621,
30674,
30726,
30777,
30827,
30877,
30926,
30975,
31023,
31070,
31117,
31163,
31209,
31253,
31298,
31341,
31384,
31426,
31468,
31509,
31549,
31589,
31628,
31666,
31704,
31741,
31778,
31813,
31849,
31883,
31917,
31950,
31983,
32015,
32046,
32076,
32106,
32136,
32164,
32192,
32219,
32246,
32272,
32297,
32322,
32346,
32369,
32392,
32414,
32435,
32456,
32476,
32495,
32514,
32532,
32550,
32566,
32582,
32598,
32612,
32626,
32640,
32652,
32665,
32676,
32687,
32697,
32706,
32715,
32723,
32730,
32737,
32743,
32748,
32753,
32757,
32760,
32763,
32765,
32766,
32767,
32767,
32766,
32765,
32763,
32760,
32757,
32753,
32748,
32743,
32737,
32730,
32723,
32715,
32706,
32697,
32687,
32676,
32665,
32652,
32640,
32626,
32612,
32598,
32582,
32566,
32550,
32532,
32514,
32495,
32476,
32456,
32435,
32414,
32392,
32369,
32346,
32322,
32297,
32272,
32246,
32219,
32192,
32164,
32136,
32106,
32076,
32046,
32015,
31983,
31950,
31917,
31883,
31849,
31813,
31778,
31741,
31704,
31666,
31628,
31589,
31549,
31509,
31468,
31426,
31384,
31341,
31298,
31253,
31209,
31163,
31117,
31070,
31023,
30975,
30926,
30877,
30827,
30777,
30726,
30674,
30621,
30568,
30515,
30460,
30406,
30350,
30294,
30237,
30180,
30122,
30063,
30004,
29944,
29884,
29823,
29761,
29699,
29636,
29572,
29508,
29443,
29378,
29312,
29246,
29179,
29111,
29043,
28974,
28904,
28834,
28764,
28692,
28621,
28548,
28475,
28402,
28327,
28253,
28177,
28101,
28025,
27948,
27870,
27792,
27713,
27634,
27554,
27474,
27393,
27311,
27229,
27146,
27063,
26979,
26895,
26810,
26725,
26639,
26552,
26465,
26378,
26290,
26201,
26112,
26022,
25932,
25841,
25749,
25658,
25565,
25472,
25379,
25285,
25190,
25095,
25000,
24904,
24807,
24710,
24613,
24515,
24416,
24317,
24218,
24118,
24017,
23916,
23815,
23713,
23610,
23507,
23404,
23300,
23196,
23091,
22985,
22880,
22773,
22667,
22559,
22452,
22344,
22235,
22126,
22017,
21907,
21796,
21686,
21574,
21463,
21350,
21238,
21125,
21011,
20898,
20783,
20668,
20553,
20438,
20322,
20205,
20089,
19971,
19854,
19736,
19617,
19498,
19379,
19260,
19140,
19019,
18898,
18777,
18656,
18534,
18411,
18289,
18165,
18042,
17918,
17794,
17669,
17544,
17419,
17294,
17168,
17041,
16915,
16788,
16660,
16532,
16404,
16276,
16147,
16018,
15889,
15759,
15629,
15499,
15368,
15237,
15106,
14974,
14842,
14710,
14578,
14445,
14312,
14178,
14045,
13911,
13776,
13642,
13507,
13372,
13237,
13101,
12965,
12829,
12693,
12556,
12419,
12282,
12144,
12007,
11869,
11730,
11592,
11453,
11315,
11175,
11036,
10896,
10757,
10617,
10476,
10336,
10195,
10054,
9913,
9772,
9631,
9489,
9347,
9205,
9063,
8920,
8778,
8635,
8492,
8349,
8205,
8062,
7918,
7775,
7631,
7486,
7342,
7198,
7053,
6908,
6764,
6619,
6473,
6328,
6183,
6037,
5892,
5746,
5600,
5454,
5308,
5162,
5015,
4869,
4722,
4576,
4429,
4282,
4135,
3988,
3841,
3694,
3547,
3400,
3252,
3105,
2957,
2810,
2662,
2515,
2367,
2219,
2071,
1923,
1776,
1628,
1480,
1332,
1184,
1036,
888,
740,
591,
443,
295,
147,
0,
-148,
-296,
-444,
-592,
-741,
-889,
-1037,
-1185,
-1333,
-1481,
-1629,
-1777,
-1924,
-2072,
-2220,
-2368,
-2516,
-2663,
-2811,
-2958,
-3106,
-3253,
-3401,
-3548,
-3695,
-3842,
-3989,
-4136,
-4283,
-4430,
-4577,
-4723,
-4870,
-5016,
-5163,
-5309,
-5455,
-5601,
-5747,
-5893,
-6038,
-6184,
-6329,
-6474,
-6620,
-6765,
-6909,
-7054,
-7199,
-7343,
-7487,
-7632,
-7776,
-7919,
-8063,
-8206,
-8350,
-8493,
-8636,
-8779,
-8921,
-9064,
-9206,
-9348,
-9490,
-9632,
-9773,
-9914,
-10055,
-10196,
-10337,
-10477,
-10618,
-10758,
-10897,
-11037,
-11176,
-11316,
-11454,
-11593,
-11731,
-11870,
-12008,
-12145,
-12283,
-12420,
-12557,
-12694,
-12830,
-12966,
-13102,
-13238,
-13373,
-13508,
-13643,
-13777,
-13912,
-14046,
-14179,
-14313,
-14446,
-14579,
-14711,
-14843,
-14975,
-15107,
-15238,
-15369,
-15500,
-15630,
-15760,
-15890,
-16019,
-16148,
-16277,
-16405,
-16533,
-16661,
-16789,
-16916,
-17042,
-17169,
-17295,
-17420,
-17545,
-17670,
-17795,
-17919,
-18043,
-18166,
-18290,
-18412,
-18535,
-18657,
-18778,
-18899,
-19020,
-19141,
-19261,
-19380,
-19499,
-19618,
-19737,
-19855,
-19972,
-20090,
-20206,
-20323,
-20439,
-20554,
-20669,
-20784,
-20899,
-21012,
-21126,
-21239,
-21351,
-21464,
-21575,
-21687,
-21797,
-21908,
-22018,
-22127,
-22236,
-22345,
-22453,
-22560,
-22668,
-22774,
-22881,
-22986,
-23092,
-23197,
-23301,
-23405,
-23508,
-23611,
-23714,
-23816,
-23917,
-24018,
-24119,
-24219,
-24318,
-24417,
-24516,
-24614,
-24711,
-24808,
-24905,
-25001,
-25096,
-25191,
-25286,
-25380,
-25473,
-25566,
-25659,
-25750,
-25842,
-25933,
-26023,
-26113,
-26202,
-26291,
-26379,
-26466,
-26553,
-26640,
-26726,
-26811,
-26896,
-26980,
-27064,
-27147,
-27230,
-27312,
-27394,
-27475,
-27555,
-27635,
-27714,
-27793,
-27871,
-27949,
-28026,
-28102,
-28178,
-28254,
-28328,
-28403,
-28476,
-28549,
-28622,
-28693,
-28765,
-28835,
-28905,
-28975,
-29044,
-29112,
-29180,
-29247,
-29313,
-29379,
-29444,
-29509,
-29573,
-29637,
-29700,
-29762,
-29824,
-29885,
-29945,
-30005,
-30064,
-30123,
-30181,
-30238,
-30295,
-30351,
-30407,
-30461,
-30516,
-30569,
-30622,
-30675,
-30727,
-30778,
-30828,
-30878,
-30927,
-30976,
-31024,
-31071,
-31118,
-31164,
-31210,
-31254,
-31299,
-31342,
-31385,
-31427,
-31469,
-31510,
-31550,
-31590,
-31629,
-31667,
-31705,
-31742,
-31779,
-31814,
-31850,
-31884,
-31918,
-31951,
-31984,
-32016,
-32047,
-32077,
-32107,
-32137,
-32165,
-32193,
-32220,
-32247,
-32273,
-32298,
-32323,
-32347,
-32370,
-32393,
-32415,
-32436,
-32457,
-32477,
-32496,
-32515,
-32533,
-32551,
-32567,
-32583,
-32599,
-32613,
-32627,
-32641,
-32653,
-32666,
-32677,
-32688,
-32698,
-32707,
-32716,
-32724,
-32731,
-32738,
-32744,
-32749,
-32754,
-32758,
-32761,
-32764,
-32766,
-32767,
-32767,
-32767,
-32767,
-32766,
-32764,
-32761,
-32758,
-32754,
-32749,
-32744,
-32738,
-32731,
-32724,
-32716,
-32707,
-32698,
-32688,
-32677,
-32666,
-32653,
-32641,
-32627,
-32613,
-32599,
-32583,
-32567,
-32551,
-32533,
-32515,
-32496,
-32477,
-32457,
-32436,
-32415,
-32393,
-32370,
-32347,
-32323,
-32298,
-32273,
-32247,
-32220,
-32193,
-32165,
-32137,
-32107,
-32077,
-32047,
-32016,
-31984,
-31951,
-31918,
-31884,
-31850,
-31814,
-31779,
-31742,
-31705,
-31667,
-31629,
-31590,
-31550,
-31510,
-31469,
-31427,
-31385,
-31342,
-31299,
-31254,
-31210,
-31164,
-31118,
-31071,
-31024,
-30976,
-30927,
-30878,
-30828,
-30778,
-30727,
-30675,
-30622,
-30569,
-30516,
-30461,
-30407,
-30351,
-30295,
-30238,
-30181,
-30123,
-30064,
-30005,
-29945,
-29885,
-29824,
-29762,
-29700,
-29637,
-29573,
-29509,
-29444,
-29379,
-29313,
-29247,
-29180,
-29112,
-29044,
-28975,
-28905,
-28835,
-28765,
-28693,
-28622,
-28549,
-28476,
-28403,
-28328,
-28254,
-28178,
-28102,
-28026,
-27949,
-27871,
-27793,
-27714,
-27635,
-27555,
-27475,
-27394,
-27312,
-27230,
-27147,
-27064,
-26980,
-26896,
-26811,
-26726,
-26640,
-26553,
-26466,
-26379,
-26291,
-26202,
-26113,
-26023,
-25933,
-25842,
-25750,
-25659,
-25566,
-25473,
-25380,
-25286,
-25191,
-25096,
-25001,
-24905,
-24808,
-24711,
-24614,
-24516,
-24417,
-24318,
-24219,
-24119,
-24018,
-23917,
-23816,
-23714,
-23611,
-23508,
-23405,
-23301,
-23197,
-23092,
-22986,
-22881,
-22774,
-22668,
-22560,
-22453,
-22345,
-22236,
-22127,
-22018,
-21908,
-21797,
-21687,
-21575,
-21464,
-21351,
-21239,
-21126,
-21012,
-20899,
-20784,
-20669,
-20554,
-20439,
-20323,
-20206,
-20090,
-19972,
-19855,
-19737,
-19618,
-19499,
-19380,
-19261,
-19141,
-19020,
-18899,
-18778,
-18657,
-18535,
-18412,
-18290,
-18166,
-18043,
-17919,
-17795,
-17670,
-17545,
-17420,
-17295,
-17169,
-17042,
-16916,
-16789,
-16661,
-16533,
-16405,
-16277,
-16148,
-16019,
-15890,
-15760,
-15630,
-15500,
-15369,
-15238,
-15107,
-14975,
-14843,
-14711,
-14579,
-14446,
-14313,
-14179,
-14046,
-13912,
-13777,
-13643,
-13508,
-13373,
-13238,
-13102,
-12966,
-12830,
-12694,
-12557,
-12420,
-12283,
-12145,
-12008,
-11870,
-11731,
-11593,
-11454,
-11316,
-11176,
-11037,
-10897,
-10758,
-10618,
-10477,
-10337,
-10196,
-10055,
-9914,
-9773,
-9632,
-9490,
-9348,
-9206,
-9064,
-8921,
-8779,
-8636,
-8493,
-8350,
-8206,
-8063,
-7919,
-7776,
-7632,
-7487,
-7343,
-7199,
-7054,
-6909,
-6765,
-6620,
-6474,
-6329,
-6184,
-6038,
-5893,
-5747,
-5601,
-5455,
-5309,
-5163,
-5016,
-4870,
-4723,
-4577,
-4430,
-4283,
-4136,
-3989,
-3842,
-3695,
-3548,
-3401,
-3253,
-3106,
-2958,
-2811,
-2663,
-2516,
-2368,
-2220,
-2072,
-1924,
-1777,
-1629,
-1481,
-1333,
-1185,
-1037,
-889,
-741,
-592,
-444,
-296,
-1481);

end sin_lut_pkg;

package body sin_lut_pkg is

---- Example 1
--  function <function_name>  (signal <signal_name> : in <type_declaration>  ) return <type_declaration> is
--    variable <variable_name>     : <type_declaration>;
--  begin
--    <variable_name> := <signal_name> xor <signal_name>;
--    return <variable_name>; 
--  end <function_name>;

---- Example 2
--  function <function_name>  (signal <signal_name> : in <type_declaration>;
--                         signal <signal_name>   : in <type_declaration>  ) return <type_declaration> is
--  begin
--    if (<signal_name> = '1') then
--      return <signal_name>;
--    else
--      return 'Z';
--    end if;
--  end <function_name>;

---- Procedure Example
--  procedure <procedure_name>  (<type_declaration> <constant_name>  : in <type_declaration>) is
--    
--  begin
--    
--  end <procedure_name>;
 
end sin_lut_pkg;
